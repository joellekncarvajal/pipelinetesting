/*
 * |-----------------------------------------------------------------------|
 * |                                                                       |
 * |   Copyright Avery Design Systems, Inc. 2010.                          |
 * |     All Rights Reserved.       Licensed Software.                     |
 * |                                                                       |
 * |                                                                       |
 * | THIS IS UNPUBLISHED PROPRIETARY SOURCE CODE OF AVERY DESIGN SYSTEMS   |
 * | The copyright notice above does not evidence any actual or intended   |
 * | publication of such source code.                                      |
 * |                                                                       |
 * |-----------------------------------------------------------------------|
 */
/*
    Test top module instantiates interface and phy modules.
*/

`timescale 1ps/1ps
import sys::*;
parameter number_of_ports = 1; //2;
parameter number_of_masters = number_of_ports;
parameter number_of_slaves = number_of_ports;


module aaxi_uvm_test_top;
   import aaxi_pkg::*;
   import aaxi_pkg_xactor::*;
   import aaxi_pkg_test::*;
   import aaxi_pll::*;
    
   import aaxi_uvm_pkg::*;
   import uvm_pkg::*;
   
   `include "uvm_macros.svh"
   
   `include "aaxi_uvm_seq_lib.svh"
   `include "my_axi_seq_lib.svh"
   
   // Normal global pings
   bit                ARESETn = 1; // AXI Reset, Deassert=H, Assert=L
   wire               ACLK;        // AXI Clock, it was generated by pll class
   reg clk;
   
   aaxi_intf     axi_if[2](ACLK, ARESETn,,,);
   
   // bus monitor/checker0
   aaxi_monitor_wrapper monitor0 (axi_if[0]);
   defparam monitor0.ID_WIDTH= AAXI_ID_WIDTH;
   defparam monitor0.BUS_DATA_WIDTH=aaxi_pkg::AAXI_DATA_WIDTH;
   defparam monitor0.USER_SUPPORT= 5'b01001;   //11111;
   
   `ifdef AVERY_AXI3
       defparam monitor0.VER= "AXI3";
       `ifdef AVERY_ASSERT_ON
        defparam monitor0.checker0.WDEPTH=4;
       `endif
   `else
       defparam monitor0.VER= "AXI4";
   `endif
       
   
   // generate Reset signal 
   initial begin
       ARESETn= 0;
       repeat(5) @(posedge ACLK);
       ARESETn= 1;
   end
   
   initial begin
       clk=0;
       forever begin
           #100 clk = ~clk;
       end
   end
   assign ACLK = clk;
   
   //SIG_AXI INTERFACE DECLARATION
   // Write master IFs
   axi_addr_inf #(
      .ID_WIDTH     (sys::axi_port_32x32x4::AXI_ID_WIDTH),
      .ADDR_WIDTH   (sys::axi_port_32x32x4::AXI_ADDR_WIDTH)
   ) axi_mstr_waddr_inf[number_of_masters-1:0](
      .clk(clk),
      .resetn(ARESETn)
   );
   axi_data_inf #(
      .ID_WIDTH     (sys::axi_port_32x32x4::AXI_ID_WIDTH),
      .DATA_WIDTH   (sys::axi_port_32x32x4::AXI_DATA_WIDTH),
      .STRB_WIDTH   (sys::axi_port_32x32x4::AXI_STRB_WIDTH)
   ) axi_mstr_wdata_inf[number_of_masters-1:0](
      .clk(clk),
      .resetn(ARESETn)
   );
   axi_resp_inf #(
      .ID_WIDTH     (sys::axi_port_32x32x4::AXI_ID_WIDTH)
   ) axi_mstr_resp_inf[number_of_masters-1:0](
      .clk(clk),
      .resetn(ARESETn)
   );

   // Read master IFs
   axi_addr_inf #(
      .ID_WIDTH     (sys::axi_port_32x32x4::AXI_ID_WIDTH),
      .ADDR_WIDTH   (sys::axi_port_32x32x4::AXI_ADDR_WIDTH)
   ) axi_mstr_raddr_inf[number_of_masters-1:0](
      .clk(clk),
      .resetn(ARESETn)
   );
   axi_data_inf #(
      .ID_WIDTH     (sys::axi_port_32x32x4::AXI_ID_WIDTH),
      .DATA_WIDTH   (sys::axi_port_32x32x4::AXI_DATA_WIDTH),
      .STRB_WIDTH   (sys::axi_port_32x32x4::AXI_STRB_WIDTH)
   ) axi_mstr_rdata_inf[number_of_masters-1:0](
      .clk(clk),
      .resetn(ARESETn)
   );

   axi_addr_inf #( 
      .ID_WIDTH     (sys::axi_port_32x32x4::AXI_ID_WIDTH),
      .ADDR_WIDTH   (sys::axi_port_32x32x4::AXI_ADDR_WIDTH)
   )axi_slv_waddr_inf[number_of_slaves-1:0](.clk(clk), .resetn(ARESETn));

   axi_data_inf #(
      .ID_WIDTH     (sys::axi_port_32x32x4::AXI_ID_WIDTH),
      .DATA_WIDTH   (sys::axi_port_32x32x4::AXI_DATA_WIDTH),
      .STRB_WIDTH   (sys::axi_port_32x32x4::AXI_STRB_WIDTH)
     ) axi_slv_wdata_inf[number_of_slaves-1:0](.clk(clk),
                                                        .resetn(ARESETn));

   axi_resp_inf #(
      .ID_WIDTH     (sys::axi_port_32x32x4::AXI_ID_WIDTH)
   ) axi_slv_resp_inf[number_of_slaves-1:0](.clk(clk),
                                                       .resetn(ARESETn));
   
   axi_addr_inf #(
      .ID_WIDTH     (sys::axi_port_32x32x4::AXI_ID_WIDTH),
      .ADDR_WIDTH   (sys::axi_port_32x32x4::AXI_ADDR_WIDTH)
   ) axi_slv_raddr_inf[number_of_slaves-1:0](.clk(clk),
                                                        .resetn(ARESETn));

   axi_data_inf #(
      .ID_WIDTH     (sys::axi_port_32x32x4::AXI_ID_WIDTH),
      .DATA_WIDTH   (sys::axi_port_32x32x4::AXI_DATA_WIDTH),
      .STRB_WIDTH   (sys::axi_port_32x32x4::AXI_STRB_WIDTH)
   ) axi_slv_rdata_inf[number_of_slaves-1:0](.clk(clk),
                                                        .resetn(ARESETn));
   genvar i;
   generate
      for (i=0; i<number_of_masters; i++) begin
         initial begin
            uvm_config_db #(sys::axi_port_32x32x4::addr_if_t)::set(null, "uvm_test_top",
                                                                   $sformatf("mstr_agent_%0d.mstr_waddr_inf", i),
                                                                   axi_mstr_waddr_inf[i]);
            uvm_config_db #(sys::axi_port_32x32x4::addr_if_t)::set(null, "uvm_test_top",
                                                                   $sformatf("mstr_agent_%0d.mstr_raddr_inf", i),
                                                                   axi_mstr_raddr_inf[i]);
            uvm_config_db #(sys::axi_port_32x32x4::data_if_t)::set(null, "uvm_test_top",
                                                                   $sformatf("mstr_agent_%0d.mstr_wdata_inf", i),
                                                                   axi_mstr_wdata_inf[i]);
            uvm_config_db #(sys::axi_port_32x32x4::data_if_t)::set(null, "uvm_test_top",
                                                                   $sformatf("mstr_agent_%0d.mstr_rdata_inf", i),
                                                                   axi_mstr_rdata_inf[i]);
            uvm_config_db #(sys::axi_port_32x32x4::resp_if_t)::set(null, "uvm_test_top",
                                                                   $sformatf("mstr_agent_%0d.mstr_resp_inf", i),
                                                                   axi_mstr_resp_inf[i]);
         end // initial begin
      end // for (i=0; i<number_of_masters; i++)
   endgenerate
   generate
      for (i=0; i<number_of_slaves; i++) begin
         initial begin
            uvm_config_db #(sys::axi_port_32x32x4::addr_if_t)::set(null, "uvm_test_top", 
                                                      $sformatf("slv_agent_%0d.slv_waddr_inf", i),
                                                      axi_slv_waddr_inf[i]);
            uvm_config_db #(sys::axi_port_32x32x4::addr_if_t)::set(null, "uvm_test_top",
                                                      $sformatf("slv_agent_%0d.slv_raddr_inf", i),
                                                      axi_slv_raddr_inf[i]);
            uvm_config_db #(sys::axi_port_32x32x4::data_if_t)::set(null, "uvm_test_top",
                                                      $sformatf("slv_agent_%0d.slv_wdata_inf", i),
                                                      axi_slv_wdata_inf[i]);
            uvm_config_db #(sys::axi_port_32x32x4::data_if_t)::set(null, "uvm_test_top",
                                                      $sformatf("slv_agent_%0d.slv_rdata_inf", i),
                                                      axi_slv_rdata_inf[i]);
            uvm_config_db #(sys::axi_port_32x32x4::resp_if_t)::set(null, "uvm_test_top",
                                                      $sformatf("slv_agent_%0d.slv_resp_inf", i),
                                                      axi_slv_resp_inf[i]);
         end // initial begin
      end // for (i=0; i<number_of_slaves; i++)
   endgenerate

   initial begin
      // AXI Configurations
      uvm_config_db #(integer)::set(null, "", "number_of_masters", number_of_masters);
      uvm_config_db #(integer)::set(null, "", "number_of_slaves", number_of_slaves);
      
      uvm_config_db #(integer)::set(null, "", "data_width_global", 32);
      uvm_config_db #(integer)::set(null, "", "address_width_global", 32);
      uvm_config_db #(integer)::set(null, "", "id_width_global", 4);
   end

   `include "sig_tests.svh"
   `include "vip_connections.svh"

   initial begin
      run_test();
   end



   
   class aaxi_uvm_test_base extends uvm_test;
       aaxi_log test_log;
   
       aaxi_uvm_testbench  tb0;
       uvm_table_printer   printer;
       aaxi_protocol_version vers;
       aaxi_cfg_info mcfg;
       aaxi_cfg_info scfg;
       bit my_slave_is_dut = 1;
   
       `uvm_component_utils( aaxi_uvm_test_base )
   
       function new( string name = "aaxi_uvm_test_base", 
   	    uvm_component parent= null, 
   `ifdef AVERY_AXI3
   	    aaxi_protocol_version vers= AAXI3
   `else
   	    aaxi_protocol_version vers= AAXI4
   `endif
   	);
   	super.new(name, parent);
   	this.vers = vers;
           test_log= new("test_log");
       endfunction : new
   
       virtual function void build_phase(uvm_phase phase); 
   	super.build_phase(phase);
   
           if($test$plusargs("MY_SLAVE_VIP")) begin
               my_slave_is_dut = 0;
               $display("MY_SLAVE_VIP plusarg found!");
           end
   
   	// Enable transaction recording for everything
   	uvm_config_int::set(this, "*", "recording_detail", UVM_FULL);
   	uvm_config_db #(aaxi_protocol_version)::set(uvm_root::get(), "*", "vers", vers);
   	$display("BENI: vers = %0s",(vers == AAXI3)?"AAXI3" : "AAXI4");
   	// ask the sequencer not to generate random sequence at the beginning
   	tb0 = aaxi_uvm_testbench::type_id::create("tb0", this);
   	uvm_config_db #(int)::set(null, "tb0.env0.master[0].sequencer.build_phase", "count", 0);
   	uvm_config_db #(int)::set(null, "tb0.env0.slave[0].sequencer.build_phase", "count", 0);
       `ifdef AVERY_PASSIVE_SLAVE
   	uvm_config_db #(int)::set(null, "tb0.env0.psv_slave[0].sequencer.build_phase", "count", 0);
       `endif
       `ifdef AVERY_PASSIVE_MASTER
   	uvm_config_db #(int)::set(null, "tb0.env0.psv_master[0].sequencer.build_phase", "count", 0);
       `endif
   
   	// set up bfm configuration
   	bfm_config_set();
   	//uvm_config_db #(aaxi_cfg_info)::set(this, "tb0.env0.master[0].driver", "cfg_info", mcfg);
   	//uvm_config_db #(aaxi_cfg_info)::set(this, "tb0.env0.slave[0].driver", "cfg_info", scfg);
   
   	uvm_config_db #(virtual aaxi_intf)::set(this, "tb0.env0.master[0].driver", "ports", aaxi_uvm_test_top.axi_if[0]);
   	uvm_config_db #(virtual aaxi_intf)::set(this, "tb0.env0.slave[0].driver", "ports", aaxi_uvm_test_top.axi_if[0]);
       `ifdef AVERY_PASSIVE_SLAVE
   	uvm_config_db #(virtual aaxi_intf)::set(this, "tb0.env0.psv_slave[0].driver", "ports", aaxi_uvm_test_top.axi_if[0]);
       `endif
       `ifdef AVERY_PASSIVE_MASTER
   	uvm_config_db #(virtual aaxi_intf)::set(this, "tb0.env0.psv_master[0].driver", "ports", aaxi_uvm_test_top.axi_if[0]);
       `endif
   	// Create a specific depth printer for printing the created topology
   	printer = new();
   	printer.knobs.depth = 4;
       endfunction : build_phase
   
       virtual function void connect_phase(uvm_phase phase);
   	super.connect_phase(phase);
           for (int i = 0; i < AAXI_INTC_MASTER_CNT; i++ ) begin
               tb0.env0.master[i].driver.cfg_info.data_bus_bytes = aaxi_pkg::AAXI_DATA_WIDTH >> 3;
               tb0.env0.master[i].driver.cfg_info.uvm_resp = 1;    
           `ifdef FOUR_OUTSTANDING
               tb0.env0.master[i].driver.cfg_info.total_outstanding_depth= 4;
               tb0.env0.master[i].driver.cfg_info.id_outstanding_depth   = 4;
           `else
               tb0.env0.master[i].driver.cfg_info.total_outstanding_depth= 1;
               tb0.env0.master[i].driver.cfg_info.id_outstanding_depth   = 1;
           `endif
           `ifdef AVERY_AXI_USER
               tb0.env0.master[i].driver.cfg_info.opt_awuser_enable= 1;
               tb0.env0.master[i].driver.cfg_info.opt_wuser_enable = 0;
               tb0.env0.master[i].driver.cfg_info.opt_buser_enable = 0;
               tb0.env0.master[i].driver.cfg_info.opt_aruser_enable= 1;
               tb0.env0.master[i].driver.cfg_info.opt_ruser_enable = 0;
           `endif
           `ifdef AVERY_PASSIVE_MASTER
               tb0.env0.psv_master[i].driver.cfg_info.data_bus_bytes = aaxi_pkg::AAXI_DATA_WIDTH >> 3;
               tb0.env0.psv_master[i].driver.cfg_info.uvm_resp = 1;
               tb0.env0.psv_master[i].driver.cfg_info.total_outstanding_depth= 1;
               tb0.env0.psv_master[i].driver.cfg_info.id_outstanding_depth   = 1;
               tb0.env0.psv_master[i].driver.cfg_info.passive_mode   = 1;
           `endif
           end
   
           // initial memory value to be 0 for data comparision on Slave BFM
           for (int i = 0; i < AAXI_INTC_SLAVE_CNT; i++ ) begin
               tb0.env0.slave[i].driver.set("mem_uninitialized_value", 0); // default memory value
               tb0.env0.slave[i].driver.cfg_info.uvm_resp = 1; // response item returned, user shall consume them, otherwise may have memory leak
               tb0.env0.slave[i].driver.cfg_info.base_address[0] = 32'h0000_0000; // memory range of address(base <=> limit)
               tb0.env0.slave[i].driver.cfg_info.limit_address[0] = 32'hFFFF_FFFF;
               tb0.env0.slave[i].driver.cfg_info.data_bus_bytes = aaxi_pkg::AAXI_DATA_WIDTH >> 3; // bytes of data_bus the device is using
               tb0.env0.slave[i].driver.add_fifo(32'habcc +i, 4); // set fifo memory address
               tb0.env0.slave[i].driver.cfg_info.total_outstanding_depth= 1;
               tb0.env0.slave[i].driver.cfg_info.id_outstanding_depth   = 1;
               tb0.env0.slave[i].driver.cfg_info.passive_mode   = my_slave_is_dut;
           `ifdef AVERY_PASSIVE_SLAVE
               tb0.env0.psv_slave[i].driver.set("mem_uninitialized_value", 0);
               tb0.env0.psv_slave[i].driver.cfg_info.uvm_resp = 1; // response item returned, user shall consume them, otherwise may have memory leak
               tb0.env0.psv_slave[i].driver.cfg_info.base_address[0] = 32'h0000_0000;
               tb0.env0.psv_slave[i].driver.cfg_info.limit_address[0] = 32'hFFFF_FFFF;
               tb0.env0.psv_slave[i].driver.cfg_info.data_bus_bytes = aaxi_pkg::AAXI_DATA_WIDTH >> 3;
               tb0.env0.psv_slave[i].driver.add_fifo(32'habcc +i, 4);
               tb0.env0.psv_slave[i].driver.cfg_info.total_outstanding_depth= 1;
               tb0.env0.psv_slave[i].driver.cfg_info.id_outstanding_depth   = 1;
               tb0.env0.psv_slave[i].driver.cfg_info.passive_mode   = 1;
           `endif
           `ifdef AVERY_AXI_USER
               tb0.env0.slave[i].driver.cfg_info.opt_awuser_enable= 1;
               tb0.env0.slave[i].driver.cfg_info.opt_wuser_enable = 0;
               tb0.env0.slave[i].driver.cfg_info.opt_buser_enable = 0;
               tb0.env0.slave[i].driver.cfg_info.opt_aruser_enable= 1;
               tb0.env0.slave[i].driver.cfg_info.opt_ruser_enable = 0;
           `endif
           end
       endfunction
   
       function void bfm_config_set();
           // move to connect_phase
       endfunction
   
       task run_phase(uvm_phase phase);
   	//uvm_test_done.set_drain_time(this, 50);
       endtask
   
       function void end_of_elaboration_phase(uvm_phase phase);
   	`uvm_info(get_type_name(),
   	    $psprintf("Printing the test topology :\n%s", this.sprint(printer)), UVM_LOW)
       endfunction : end_of_elaboration_phase
   
       virtual function void report_phase(uvm_phase phase);
           uvm_report_server rpt = uvm_report_server::get_server();
           int  cnt1 = rpt.get_severity_count(UVM_ERROR);
           int  cnt2 = rpt.get_severity_count(UVM_FATAL);
           
           super.report_phase(phase);
   
           test_log.merge_coverage(tb0.env0.master[0].driver.log);
           test_log.merge_coverage(tb0.env0.slave[0].driver.log);
   
           // print out assertion coverage
           test_log.coverage_rpt();
   
           if (cnt1 || cnt2)                                                                                                                                                                     
               `uvm_info(get_type_name(),
                   $psprintf("Test failed due to UVM_ERROR=%0d and UVM_FATAL=%0d", cnt1, cnt2), UVM_LOW);
       endfunction : report_phase
   
   endclass: aaxi_uvm_test_base
   
   
   /*************************************************/
   /******************uvm tests *********************/
   /*************************************************/
   `include "my_axi_base_test.sv"
   `include "aaxi_uvm_example_tests.svh"
   `include "my_testlist.sv"
   
   final begin
   $display("%0t: BENI_FINAL", $time);
   end
   
//   initial begin
//   //DUMP_WAVEFORM
//   `ifdef AAXI_DUMP_VCD
//       $dumpfile("aaxi_top.vcd");
//       $dumpvars(0, aaxi_uvm_test_top);
//       $dumpon;
//       `ifdef AVERY_MS
//           `ifdef AVERY_AXI4_STREAM
//   	    $dumpvars(0, aaxi_uvm_test_top.portstream);
//           `endif
//       `endif
//   `endif
//   
//   `ifdef AAXI_DUMP_VPD
//       $vcdplusfile("aaxi_top.vpd");
//       $vcdpluson(0, aaxi_uvm_test_top);
//   `endif
//   
//   `ifdef AAXI_DUMP_FSDB
//       $fsdbDumpfile("aaxi_uvm_test_top.fsdb");
//       $fsdbDumpvars(0, aaxi_uvm_test_top, "+all");
//       $fsdbDumpon;
//   `endif
//   end
//   
//   initial begin
//     $display("BENI - AXI_ALIGN_ADDR = %0d",`AXI_ALIGN_ADDR);
//     $shm_open("waves.shm"); $shm_probe("AS");
//   end


endmodule
