`define AXI_ADDR_WIDTH 32
`define AXI_DATA_WIDTH 32
`define AXI_USER_WIDTH 1
`define AXI_ID_WIDTH 4
`define AXI_STRB_WIDTH `AXI_DATA_WIDTH/8
`define AXI_ALIGN_ADDR $clog2(`AXI_DATA_WIDTH/8)

`define AAXI_MAX_AWUSER_WIDTH `AXI_USER_WIDTH
`define AAXI_MAX_ARUSER_WIDTH `AXI_USER_WIDTH
//`define AAXI_INTC_SLAVE_CNT 0
