/*
   ######################################################################################
 *      Signature IP Corporation Confidential and Proprietary Information               #
 *      Copyright 2022 Signature IP Corporation                                         #
 *      All Rights Reserved.                                                            #
 *      This is UNPUBLISHED PROPRIETARY SOURCE CODE OF Signature IP Corporation         #
 *      The copyright notice above does not evidence any actual or intended publication #
 *      of such source code.                                                            #
 * ######################################################################################

*/
package sig_axi_pkg;
   
   import uvm_pkg::*;
   `include "uvm_macros.svh"
   import axi_pkg::*;

   `include "sig_axi_env.sv"   
   
endpackage // sig_axi_pkg
