/*
   ######################################################################################
 *      Signature IP Corporation Confidential and Proprietary Information               #
 *      Copyright 2022 Signature IP Corporation                                         #
 *      All Rights Reserved.                                                            #
 *      This is UNPUBLISHED PROPRIETARY SOURCE CODE OF Signature IP Corporation         #
 *      The copyright notice above does not evidence any actual or intended publication #
 *      of such source code.                                                            #
 * ######################################################################################

*/
`ifndef axi_driver__sv
 `define axi_driver__sv
class axi_addr_driver #(type T=axi_params)extends uvm_driver#(axi_addr_item#(
    .AXI_ID_WIDTH    (T::AXI_ID_WIDTH),
    .AXI_ADDR_WIDTH  (T::AXI_ADDR_WIDTH),
    .AXI_LEN_WIDTH   (T::AXI_LEN_WIDTH),
    .AXI_SIZE_WIDTH  (T::AXI_SIZE_WIDTH),
    .AXI_BURST_WIDTH (T::AXI_BURST_WIDTH),
    .AXI_LOCK_WIDTH  (T::AXI_LOCK_WIDTH),
    .AXI_CACHE_WIDTH (T::AXI_CACHE_WIDTH),
    .AXI_PROT_WIDTH  (T::AXI_PROT_WIDTH),
    .AXI_QOS_WIDTH   (T::AXI_QOS_WIDTH),
    .AXI_REGION_WIDTH(T::AXI_REGION_WIDTH),
    .AXI_USER_WIDTH  (T::AXI_USER_WIDTH)
));

   `uvm_component_param_utils(axi_addr_driver#(T))

   //typedef T::axi_addr_item_t axi_addr_item_type;
   //typedef T::addr_if_t addr_if_type;
   typedef axi_addr_item # (
     .AXI_ID_WIDTH     (T::AXI_ID_WIDTH), 
     .AXI_ADDR_WIDTH   (T::AXI_ADDR_WIDTH),
     .AXI_LEN_WIDTH    (T::AXI_LEN_WIDTH),
     .AXI_SIZE_WIDTH   (T::AXI_SIZE_WIDTH),
     .AXI_BURST_WIDTH  (T::AXI_BURST_WIDTH),
     .AXI_LOCK_WIDTH   (T::AXI_LOCK_WIDTH),
     .AXI_CACHE_WIDTH  (T::AXI_CACHE_WIDTH),
     .AXI_PROT_WIDTH   (T::AXI_PROT_WIDTH),
     .AXI_QOS_WIDTH    (T::AXI_QOS_WIDTH),
     .AXI_REGION_WIDTH (T::AXI_REGION_WIDTH),
     .AXI_USER_WIDTH   (T::AXI_USER_WIDTH)
   ) axi_addr_item_type;
  typedef virtual axi_addr_inf #( 
    .ID_WIDTH     (T::AXI_ID_WIDTH),
    .ADDR_WIDTH   (T::AXI_ADDR_WIDTH),
    .LEN_WIDTH    (T::AXI_LEN_WIDTH),
    .SIZE_WIDTH   (T::AXI_SIZE_WIDTH),
    .BURST_WIDTH  (T::AXI_BURST_WIDTH),
    .LOCK_WIDTH   (T::AXI_LOCK_WIDTH),
    .CACHE_WIDTH  (T::AXI_CACHE_WIDTH),
    .PROT_WIDTH   (T::AXI_PROT_WIDTH),
    .QOS_WIDTH    (T::AXI_QOS_WIDTH),
    .REGION_WIDTH (T::AXI_REGION_WIDTH),
    .USER_WIDTH   (T::AXI_USER_WIDTH),
    .GPIO_WIDTH   (T::AXI_GPIO_WIDTH)
  ) addr_if_type;

   addr_if_type addr_if;
   OpType   rwType;
   bit req_ongoing; 
   bit do_sw_reset = 0;
   axi_port_cfg cfg;

   function new(string name="axi_addr_driver", uvm_component parent=null);
      super.new(name, parent);
   endfunction // new

   `protect //begin protected region
   function void print_params();
      $display("%0s params:", get_full_name());
      $display("AXI_ID_WIDTH     = %0d",    T::AXI_ID_WIDTH);
      $display("AXI_ADDR_WIDTH   = %0d",  T::AXI_ADDR_WIDTH);
      $display("AXI_LEN_WIDTH    = %0d",   T::AXI_LEN_WIDTH);
      $display("AXI_SIZE_WIDTH   = %0d",  T::AXI_SIZE_WIDTH);
      $display("AXI_BURST_WIDTH  = %0d", T::AXI_BURST_WIDTH);
      $display("AXI_LOCK_WIDTH   = %0d",  T::AXI_LOCK_WIDTH);
      $display("AXI_CACHE_WIDTH  = %0d", T::AXI_CACHE_WIDTH);
      $display("AXI_PROT_WIDTH   = %0d",  T::AXI_PROT_WIDTH);
      $display("AXI_QOS_WIDTH    = %0d",   T::AXI_QOS_WIDTH);
      $display("AXI_REGION_WIDTH = %0d",T::AXI_REGION_WIDTH);
      $display("AXI_USER_WIDTH   = %0d",  T::AXI_USER_WIDTH);
      $display("AXI_WR_ID_WIDTH  = %0d",    T::AXI_WR_ID_WIDTH);
      $display("AXI_RD_ID_WIDTH  = %0d",    T::AXI_RD_ID_WIDTH);
   endfunction

   virtual function void build_phase(uvm_phase phase);
      super.build_phase(phase);
      //print_params();
   endfunction // build_phase
   
   virtual function void connect_phase(uvm_phase phase);
      super.connect_phase(phase);
   endfunction // connect_phase
   
   task reset_phase(uvm_phase phase);
      //phase.raise_objection(this);
      //super.reset_phase(phase);
      //addr_if.src_drv_cb.AxVALID <= 'h0;
      //addr_if.src_drv_cb.AxID    <= 'h0;
      //addr_if.src_drv_cb.AxADDR  <= 'h0;
      //addr_if.src_drv_cb.AxLEN   <= 'h0;
      //addr_if.src_drv_cb.AxSIZE  <= 'h0;
      //addr_if.src_drv_cb.AxBURST <= 'h0;
      //addr_if.src_drv_cb.AxLOCK  <= 'h0;
      //addr_if.src_drv_cb.AxCACHE <= 'h0;
      //addr_if.src_drv_cb.AxPROT  <= 'h0;
      //addr_if.src_drv_cb.AxQOS   <= 'h0;
      //addr_if.src_drv_cb.AxREGION<= 'h0;
      //addr_if.src_drv_cb.AxUSER  <= 'h0;
      //addr_if.src_drv_cb.AxGPIO  <= 'h0;
      ////`uvm_info(get_name(), "Waiting for resetn deassertion...", UVM_NONE)      
      ////wait(addr_if.src_drv_cb.resetn == 1'b1);
      ////repeat(10) @(addr_if.src_drv_cb);
      ////`uvm_info(get_name(), "AXI_RESET_N deasserts", UVM_LOW)
      //phase.drop_objection(this);
   endtask // reset_phase

   task reset_handler();
      //$display("%0t: %0s reset_handler", $time, get_full_name());
      while (addr_if.src_drv_cb.resetn === 1'b1) begin
         @(addr_if.src_drv_cb);
      end
      addr_if.src_drv_cb.AxVALID <= 'h0;
      addr_if.src_drv_cb.AxID    <= 'h0;
      addr_if.src_drv_cb.AxADDR  <= 'h0;
      addr_if.src_drv_cb.AxLEN   <= 'h0;
      addr_if.src_drv_cb.AxSIZE  <= 'h0;
      addr_if.src_drv_cb.AxBURST <= 'h0;
      addr_if.src_drv_cb.AxLOCK  <= 'h0;
      addr_if.src_drv_cb.AxCACHE <= 'h0;
      addr_if.src_drv_cb.AxPROT  <= 'h0;
      addr_if.src_drv_cb.AxQOS   <= 'h0;
      addr_if.src_drv_cb.AxREGION<= 'h0;
      addr_if.src_drv_cb.AxUSER  <= 'h0;
      addr_if.src_drv_cb.AxGPIO  <= 'h0;
      if (req_ongoing == 1) begin
         seq_item_port.item_done(req);
         req_ongoing = 0;
      end
   endtask

   task sw_reset_seq();
      while (do_sw_reset == 0) begin
         @(addr_if.src_drv_cb);
      end
      addr_if.src_drv_cb.AxVALID <= 'h0;
      addr_if.src_drv_cb.AxID    <= 'h0;
      addr_if.src_drv_cb.AxADDR  <= 'h0;
      addr_if.src_drv_cb.AxLEN   <= 'h0;
      addr_if.src_drv_cb.AxSIZE  <= 'h0;
      addr_if.src_drv_cb.AxBURST <= 'h0;
      addr_if.src_drv_cb.AxLOCK  <= 'h0;
      addr_if.src_drv_cb.AxCACHE <= 'h0;
      addr_if.src_drv_cb.AxPROT  <= 'h0;
      addr_if.src_drv_cb.AxQOS   <= 'h0;
      addr_if.src_drv_cb.AxREGION<= 'h0;
      addr_if.src_drv_cb.AxUSER  <= 'h0;
      addr_if.src_drv_cb.AxGPIO  <= 'h0;
      if (req_ongoing == 1) begin
         seq_item_port.item_done(req);
         req_ongoing = 0;
      end
      //do_sw_reset = 0;
   endtask

   task drain_sqr();
      axi_addr_item_type tr;

      if (req_ongoing == 1) begin
         seq_item_port.item_done();
         req_ongoing = 0;
      end
      do begin
         seq_item_port.try_next_item(tr);
         if ((tr != null)) seq_item_port.item_done();
      end while (tr != null);      
   endtask

   task drive_rand_value();
      axi_addr_item_type rand_addr;
      rand_addr = axi_addr_item_type::type_id::create("rand_addr", this);
      rand_addr.randomize();  
      addr_if.src_drv_cb.AxVALID <= 1'b0;
      addr_if.src_drv_cb.AxID    <= rand_addr.id;
      addr_if.src_drv_cb.AxADDR  <= rand_addr.addr;
      addr_if.src_drv_cb.AxLEN   <= rand_addr.len;
      addr_if.src_drv_cb.AxSIZE  <= rand_addr.size;
      addr_if.src_drv_cb.AxBURST <= rand_addr.burst;
      addr_if.src_drv_cb.AxLOCK  <= rand_addr.lock;
      addr_if.src_drv_cb.AxCACHE <= rand_addr.cache;
      addr_if.src_drv_cb.AxPROT  <= rand_addr.prot;
      addr_if.src_drv_cb.AxQOS   <= rand_addr.qos;
      addr_if.src_drv_cb.AxREGION<= rand_addr.region;
      addr_if.src_drv_cb.AxUSER  <= rand_addr.user;
      addr_if.src_drv_cb.AxGPIO  <= rand_addr.gpio;
   endtask

   task drive_if();
      axi_addr_item_type tr;
      int delay_cnt = 0;
      bit[T::AXI_ID_WIDTH-1:0] actual_id;

      req_ongoing = 0;
      while(addr_if.src_drv_cb.resetn !== 1'b1) begin
         @(addr_if.src_drv_cb);
      end
      forever begin
         //seq_item_port.get_next_item(tr);
         seq_item_port.try_next_item(tr);
         while (tr == null) begin
            if (cfg.en_rand_while_not_valid == 1'b1) drive_rand_value();
            @(addr_if.src_drv_cb);
            seq_item_port.try_next_item(tr);
         end
         tr.rwType = rwType;
         //CONFIGURABLE WR/RD ID WIDTHS
         actual_id = '0;
         if (rwType == WRITE) begin
            if (T::AXI_ID_WIDTH > T::AXI_WR_ID_WIDTH) begin
               actual_id[T::AXI_WR_ID_WIDTH-1:0] = tr.id[T::AXI_WR_ID_WIDTH-1:0];
            end else begin
               actual_id = tr.id;
            end
         end else if (rwType == READ) begin
            if (T::AXI_ID_WIDTH > T::AXI_RD_ID_WIDTH) begin
               actual_id[T::AXI_RD_ID_WIDTH-1:0] = tr.id[T::AXI_RD_ID_WIDTH-1:0];
            end else begin
               actual_id = tr.id;
            end
         end
         //CONFIGURABLE WR/RD ID WIDTHS
         `uvm_info(get_full_name(), $sformatf("Starting transaction: %s", tr.sprint()), UVM_DEBUG)
         req_ongoing = 1;
         //insert delay handling here
         repeat (tr.delay) @(addr_if.src_drv_cb);
         delay_cnt = 0; //Used for timeout
         addr_if.src_drv_cb.AxVALID <= 1'b1;
         addr_if.src_drv_cb.AxID    <= actual_id; //tr.id; //CONFIGURABLE WR/RD ID WIDTHS
         addr_if.src_drv_cb.AxADDR  <= tr.addr;
         addr_if.src_drv_cb.AxLEN   <= tr.len;
         addr_if.src_drv_cb.AxSIZE  <= tr.size;
         addr_if.src_drv_cb.AxBURST <= tr.burst;
         addr_if.src_drv_cb.AxLOCK  <= tr.lock;
         addr_if.src_drv_cb.AxCACHE <= tr.cache;
         addr_if.src_drv_cb.AxPROT  <= tr.prot;
         addr_if.src_drv_cb.AxQOS   <= tr.qos;
         addr_if.src_drv_cb.AxREGION<= tr.region;
         addr_if.src_drv_cb.AxUSER  <= tr.user;
	 addr_if.src_drv_cb.AxGPIO  <= tr.gpio;
         @(addr_if.src_drv_cb);
         while(addr_if.src_drv_cb.AxREADY == 0 && delay_cnt <= T::READY_TIMEOUT) begin
            @(addr_if.src_drv_cb);
            delay_cnt++;
         end
         if (delay_cnt > T::READY_TIMEOUT) begin
            `uvm_fatal("READY_TIMEOUT",$sformatf("Timeout while waiting for ready signal to assert. %0d cycles passed while waiting for ready.", delay_cnt));
         end
         addr_if.src_drv_cb.AxVALID <= 1'b0;
         req_ongoing = 0;
         seq_item_port.item_done();
      end // forever
   endtask

   task run_phase(uvm_phase phase);
      @(addr_if.src_drv_cb);
      forever begin
         fork
            begin
               fork
                  reset_handler();
                  drive_if();
                  sw_reset_seq();
               join_any
            end
         join
         disable fork;
         while (addr_if.src_drv_cb.resetn !== 1 || do_sw_reset == 1) begin
            @(addr_if.src_drv_cb);
         end //while
      end //forever
   endtask

   `endprotect //end protected region
endclass // axi_addr_driver

class axi_data_driver #(type T=axi_params) extends uvm_driver#(axi_data_item#(
    .AXI_ID_WIDTH  (T::AXI_ID_WIDTH),
    .AXI_DATA_WIDTH(T::AXI_DATA_WIDTH),
    .AXI_STRB_WIDTH(T::AXI_STRB_WIDTH),
    .AXI_RESP_WIDTH(T::AXI_RESP_WIDTH),
    .AXI_USER_WIDTH  (T::AXI_USER_WIDTH)
));


   `uvm_component_param_utils(axi_data_driver#(T))
   //typedef T::axi_data_item_t axi_data_item_type;
   //typedef T::data_if_t data_if_type;
   typedef axi_data_item#(
     .AXI_ID_WIDTH(T::AXI_ID_WIDTH),
     .AXI_DATA_WIDTH(T::AXI_DATA_WIDTH),
     .AXI_STRB_WIDTH(T::AXI_STRB_WIDTH),
     .AXI_RESP_WIDTH(T::AXI_RESP_WIDTH),
     .AXI_USER_WIDTH(T::AXI_USER_WIDTH)
   ) axi_data_item_type;
  typedef virtual axi_data_inf #(
    .ID_WIDTH     (T::AXI_ID_WIDTH),
    .DATA_WIDTH   (T::AXI_DATA_WIDTH), 
    .STRB_WIDTH   (T::AXI_STRB_WIDTH),
    .USER_WIDTH   (T::AXI_USER_WIDTH),
    .RESP_WIDTH   (T::AXI_RESP_WIDTH)
  ) data_if_type;

   OpType   rwType;
   data_if_type data_if;
   bit req_ongoing;
   axi_port_cfg cfg;

   function new(string name="axi_data_driver", uvm_component parent=null);
      super.new(name, parent);
   endfunction // new

   `protect //begin protected region
   function void print_params();
      $display("%0s params:", get_full_name());
      $display("AXI_ID_WIDTH   = %0d",    T::AXI_ID_WIDTH);
      $display("AXI_DATA_WIDTH = %0d",T::AXI_DATA_WIDTH);
      $display("AXI_STRB_WIDTH = %0d",T::AXI_STRB_WIDTH);
      $display("AXI_RESP_WIDTH = %0d",T::AXI_RESP_WIDTH);
   endfunction

   virtual function void build_phase(uvm_phase phase);
      super.build_phase(phase);
      //print_params();
   endfunction // build_phase
   
   virtual function void connect_phase(uvm_phase phase);
      super.connect_phase(phase);
   endfunction // connect_phase
   
   task drive_rand_value();
      axi_data_item_type rand_data;
      rand_data = axi_data_item_type::type_id::create("rand_data", this);
      rand_data.randomize() with {
         data.size() == 1;
         strb.size() == 1;
         user.size() == 1;
         resp.size() == 1;
         delay.size() == 1;
      };
      data_if.src_drv_cb.xVALID <= 'h0;
      data_if.src_drv_cb.xID    <= rand_data.id;
      data_if.src_drv_cb.xDATA  <= rand_data.data[0];
      data_if.src_drv_cb.xLAST  <= ^(rand_data.data[0]);
      if (rwType == READ) begin
         data_if.src_drv_cb.xRESP  <= rand_data.resp[0];
      end else if (rwType == WRITE) begin
         data_if.src_drv_cb.xSTRB  <= rand_data.strb[0];
      end
      data_if.src_drv_cb.xUSER  <= rand_data.user[0];
   endtask

   task reset_phase(uvm_phase phase);
      //phase.raise_objection(this);
      //super.reset_phase(phase);
      //data_if.src_drv_cb.xVALID <= 'h0;
      //data_if.src_drv_cb.xID    <= 'h0;
      //data_if.src_drv_cb.xDATA  <= 'h0;
      //data_if.src_drv_cb.xSTRB  <= 'h0;
      //data_if.src_drv_cb.xLAST  <= 'h0;
      //data_if.src_drv_cb.xRESP  <= 'h0;
      //data_if.src_drv_cb.xUSER  <= 'h0;
      ////wait(data_if.src_drv_cb.resetn == 1'b1);
      ////repeat(10) @(posedge data_if.clk);
      ////`uvm_info(get_name(), "AXI_RESET_N deasserts", UVM_LOW)
      //phase.drop_objection(this);
   endtask // reset_phase

   task reset_handler();
      while (data_if.src_drv_cb.resetn === 1'b1  
            //&& ((cfg.rdata_ch_is_unresponsive == '0 && rwType == READ) || (cfg.wdata_ch_is_unresponsive == '0 && rwType == WRITE))
      ) begin
         @(data_if.src_drv_cb);
      end
      data_if.src_drv_cb.xVALID <= 'h0;
      data_if.src_drv_cb.xID    <= 'h0;
      data_if.src_drv_cb.xDATA  <= 'h0;
      data_if.src_drv_cb.xSTRB  <= 'h0;
      data_if.src_drv_cb.xLAST  <= 'h0;
      data_if.src_drv_cb.xRESP  <= 'h0;
      data_if.src_drv_cb.xUSER  <= 'h0;
      if (req_ongoing == 1) begin
         seq_item_port.item_done(req);
      end
   endtask

   task drive_if();
      axi_data_item_type tr;
      int unsigned delay_cnt = 0, data_cnt;
      bit[T::AXI_ID_WIDTH-1:0] actual_id;

      req_ongoing = 0;
      while(data_if.src_drv_cb.resetn !== 1'b1) begin
         @(data_if.src_drv_cb);
      end
      forever begin
         //seq_item_port.get_next_item(tr);
         //while ((cfg.rdata_ch_is_unresponsive == 1'b1 && rwType == READ) || (cfg.wdata_ch_is_unresponsive == 1'b1 && rwType == WRITE)) begin
         //   @(data_if.src_drv_cb);
         //end
         while (cfg.pause_rdata_ch == 1'b1 && rwType == READ) begin
            @(data_if.src_drv_cb);
         end 
         seq_item_port.try_next_item(tr);
         while (tr == null) begin
            if (cfg.en_rand_while_not_valid == 1'b1) drive_rand_value();
            @(data_if.src_drv_cb);
            seq_item_port.try_next_item(tr);
         end
         tr.rwType = rwType;
         //CONFIGURABLE WR/RD ID WIDTHS
         actual_id = '0;
         if (rwType == WRITE) begin
            if (T::AXI_ID_WIDTH > T::AXI_WR_ID_WIDTH) begin
               actual_id[T::AXI_WR_ID_WIDTH-1:0] = tr.id[T::AXI_WR_ID_WIDTH-1:0];
            end else begin
               actual_id = tr.id;
            end
         end else if (rwType == READ) begin
            if (T::AXI_ID_WIDTH > T::AXI_RD_ID_WIDTH) begin
               actual_id[T::AXI_RD_ID_WIDTH-1:0] = tr.id[T::AXI_RD_ID_WIDTH-1:0];
            end else begin
               actual_id = tr.id;
            end
         end
         //CONFIGURABLE WR/RD ID WIDTHS

         `uvm_info(get_full_name(), $sformatf("Starting transaction: %s", tr.sprint()), UVM_DEBUG)
         req_ongoing = 1;
         delay_cnt = 0; //Used for timeout
         //Driving logic
         data_cnt = 0;
         while (data_cnt != tr.data_len &&
               ((cfg.rdata_ch_is_unresponsive == 1'b0 && rwType == READ) || (cfg.wdata_ch_is_unresponsive == 1'b0 && rwType == WRITE))
         ) begin
            //insert delay per beat
            repeat (tr.delay[data_cnt]) @(data_if.src_drv_cb);
            data_if.src_drv_cb.xVALID <= 1'b1;
            data_if.src_drv_cb.xID <= actual_id; //tr.id; //[data_cnt];  //May need to use array for ID to support interleave
            data_if.src_drv_cb.xDATA <= tr.data[data_cnt];
            if (data_cnt == tr.data_len-1 && tr.not_last == 0) begin
               data_if.src_drv_cb.xLAST <= 1'b1;
            end else begin
               data_if.src_drv_cb.xLAST <= 1'b0;
            end
            if (tr.rwType == READ) begin
               data_if.src_drv_cb.xRESP <= tr.resp[data_cnt];
            end else begin
               data_if.src_drv_cb.xSTRB <= tr.strb[data_cnt];
            end
            data_if.src_drv_cb.xUSER <= tr.user[data_cnt];
            @(data_if.src_drv_cb);
            data_cnt++;
            while (data_if.src_drv_cb.xREADY == 1'b0 && delay_cnt <= T::READY_TIMEOUT) begin
               @(data_if.src_drv_cb);
               delay_cnt++;
            end
            if (delay_cnt > T::READY_TIMEOUT) begin
            `uvm_fatal("READY_TIMEOUT",$sformatf("Timeout while waiting for ready signal to assert. %0d cycles passed while waiting for ready.", delay_cnt));
            end //if
            data_if.src_drv_cb.xVALID <= 1'b0;
            delay_cnt=0; //reset timeout counter
         end //while
         req_ongoing = 0;
         seq_item_port.item_done();
      end
   endtask

   task run_phase(uvm_phase phase);
      @(data_if.src_drv_cb);
      forever begin
         fork
            begin
               fork
                  reset_handler();
                  drive_if();
               join_any
            end
         join
         disable fork;
         while (data_if.src_drv_cb.resetn !== 1  
               //|| ((cfg.rdata_ch_is_unresponsive == 1'b1 && rwType == READ) || (cfg.wdata_ch_is_unresponsive == 1'b1 && rwType == WRITE))
         ) begin
            @(data_if.src_drv_cb);
         end //while
      end //forever
   endtask

   `endprotect //end protected region
endclass // axi_addr_driver

class axi_resp_driver #(type T=axi_params) extends uvm_driver#(axi_resp_item#(
    .AXI_ID_WIDTH  (T::AXI_ID_WIDTH),
    .AXI_RESP_WIDTH(T::AXI_RESP_WIDTH),
    .AXI_USER_WIDTH(T::AXI_USER_WIDTH)
));

   `uvm_component_param_utils(axi_resp_driver#(T))
   //typedef T::axi_resp_item_t axi_resp_item_type;
   //typedef T::resp_if_t resp_if_type;
   typedef axi_resp_item #(
     .AXI_ID_WIDTH (T::AXI_ID_WIDTH),
     .AXI_RESP_WIDTH (T::AXI_RESP_WIDTH),
     .AXI_USER_WIDTH (T::AXI_USER_WIDTH)
   ) axi_resp_item_type;
  typedef virtual axi_resp_inf #(
    .ID_WIDTH     (T::AXI_ID_WIDTH),
    .RESP_WIDTH   (T::AXI_RESP_WIDTH),
    .USER_WIDTH   (T::AXI_USER_WIDTH)
  ) resp_if_type;

   resp_if_type resp_if;
   OpType rwType;
   bit req_ongoing;
   axi_port_cfg cfg;

   function new(string name="axi_resp_driver", uvm_component parent=null);
      super.new(name, parent);
   endfunction // new

   `protect //begin protected region
   function void print_params();
      $display("%0s params:", get_full_name());
      $display("AXI_ID_WIDTH   = %0d",    T::AXI_ID_WIDTH);
      $display("AXI_RESP_WIDTH = %0d",T::AXI_RESP_WIDTH);
   endfunction

   virtual function void build_phase(uvm_phase phase);
      super.build_phase(phase);
      //print_params();
   endfunction // build_phase
   
   virtual function void connect_phase(uvm_phase phase);
      super.connect_phase(phase);
   endfunction // connect_phase
   
   task reset_phase(uvm_phase phase);
   endtask // reset_phase

   task drive_rand_value();
      axi_resp_item_type rand_resp;
      rand_resp = axi_resp_item_type::type_id::create("rand_resp", this);
      rand_resp.randomize();
      resp_if.src_drv_cb.BVALID <= 'h0;
      resp_if.src_drv_cb.BID    <= rand_resp.id;
      resp_if.src_drv_cb.BRESP  <= rand_resp.resp;
      resp_if.src_drv_cb.BUSER  <= rand_resp.user;
   endtask

   task reset_handler();
      while (resp_if.src_drv_cb.resetn === 1'b1) begin
         @(resp_if.src_drv_cb);
      end
      resp_if.src_drv_cb.BVALID <= 'h0;
      resp_if.src_drv_cb.BID    <= 'h0;
      resp_if.src_drv_cb.BRESP  <= 'h0;
      resp_if.src_drv_cb.BUSER  <= 'h0;
      if (req_ongoing == 1) begin
         seq_item_port.item_done(req);
      end
   endtask

   task drive_if();
      axi_resp_item_type tr;
      int unsigned delay_cnt = 0;
      bit[T::AXI_ID_WIDTH-1:0] actual_id;

      req_ongoing = 0;
      while(resp_if.src_drv_cb.resetn !== 1'b1) begin
         @(resp_if.src_drv_cb);
      end
      forever begin
         //seq_item_port.get_next_item(tr);
         while (cfg.pause_bresp_ch == 1'b1) begin
            @(resp_if.src_drv_cb);
         end
         seq_item_port.try_next_item(tr);
         while (tr == null) begin
            if (cfg.en_rand_while_not_valid == 1'b1) drive_rand_value();
            @(resp_if.src_drv_cb);
            seq_item_port.try_next_item(tr);
         end
         tr.rwType = rwType;
         //CONFIGURABLE WR/RD ID WIDTHS
         actual_id = '0;
         //$display("ACTUAL_ID_DBG: AXI_ID_WIDTH=%0d, AXI_WR_ID_WIDTH=%0d", T::AXI_ID_WIDTH, T::AXI_WR_ID_WIDTH);
         if (T::AXI_ID_WIDTH > T::AXI_WR_ID_WIDTH) begin
            actual_id[T::AXI_WR_ID_WIDTH-1:0] = tr.id[T::AXI_WR_ID_WIDTH-1:0];
         end else begin
            actual_id = tr.id;
         end
         //CONFIGURABLE WR/RD ID WIDTHS

         `uvm_info(get_full_name(), $sformatf("Starting transaction: %s", tr.sprint()), UVM_DEBUG)
         req_ongoing = 1;

      if (cfg.bresp_ch_is_unresponsive == 0) begin   
         //insert delay handling here
         repeat (tr.delay) @(resp_if.src_drv_cb);
         delay_cnt = 0; //Used for timeout

         //Driving logic
         resp_if.src_drv_cb.BVALID <= 1'b1;
         resp_if.src_drv_cb.BID    <= actual_id; //tr.id;
         resp_if.src_drv_cb.BRESP  <= tr.resp; //[0];
         resp_if.src_drv_cb.BUSER  <= tr.user;
         @(resp_if.src_drv_cb);
         while (resp_if.src_drv_cb.BREADY == 0 && delay_cnt <= T::READY_TIMEOUT) begin
            @(resp_if.src_drv_cb);
            delay_cnt++;
         end
         if (delay_cnt > T::READY_TIMEOUT) begin
            `uvm_fatal("READY_TIMEOUT",$sformatf("Timeout while waiting for ready signal to assert. %0d cycles passed while waiting for ready.", delay_cnt));
         end //if
      end
         resp_if.src_drv_cb.BVALID <= 1'b0;
         req_ongoing = 0;
         seq_item_port.item_done();
      end //forever
   endtask


   task run_phase(uvm_phase phase);
      @(resp_if.src_drv_cb);
      forever begin
         fork
            begin
               fork
                  reset_handler();
                  drive_if();
               join_any
            end
         join
         disable fork;
         while (resp_if.src_drv_cb.resetn !== 1) begin
            @(resp_if.src_drv_cb);
         end //while
      end //forever
   endtask // run_phase

   `endprotect //end protected region
endclass // axi_resp_driver

class axi_ready_driver#(type T=axi_params) extends uvm_component;
   `uvm_component_param_utils(axi_ready_driver#(T))

   //typedef T::addr_if_t addr_if_type;
   //typedef T::data_if_t data_if_type;
   //typedef T::resp_if_t resp_if_type;
  typedef virtual axi_addr_inf #( 
    .ID_WIDTH     (T::AXI_ID_WIDTH),
    .ADDR_WIDTH   (T::AXI_ADDR_WIDTH),
    .LEN_WIDTH    (T::AXI_LEN_WIDTH),
    .SIZE_WIDTH   (T::AXI_SIZE_WIDTH),
    .BURST_WIDTH  (T::AXI_BURST_WIDTH),
    .LOCK_WIDTH   (T::AXI_LOCK_WIDTH),
    .CACHE_WIDTH  (T::AXI_CACHE_WIDTH),
    .PROT_WIDTH   (T::AXI_PROT_WIDTH),
    .QOS_WIDTH    (T::AXI_QOS_WIDTH),
    .REGION_WIDTH (T::AXI_REGION_WIDTH),
    .USER_WIDTH   (T::AXI_USER_WIDTH),
    .GPIO_WIDTH   (T::AXI_GPIO_WIDTH)
  ) addr_if_type;

  typedef virtual axi_data_inf #(
    .ID_WIDTH     (T::AXI_ID_WIDTH),
    .DATA_WIDTH   (T::AXI_DATA_WIDTH), 
    .STRB_WIDTH   (T::AXI_STRB_WIDTH),
    .USER_WIDTH   (T::AXI_USER_WIDTH),
    .RESP_WIDTH   (T::AXI_RESP_WIDTH)
  ) data_if_type;

  typedef virtual axi_resp_inf #(
    .ID_WIDTH     (T::AXI_ID_WIDTH),
    .RESP_WIDTH   (T::AXI_RESP_WIDTH),
    .USER_WIDTH   (T::AXI_USER_WIDTH)
  ) resp_if_type;

   ChType channelType;
   OpType direction;
   int min_ready_delay=0, max_ready_delay=0;
   int ready_high_cycles;
   addr_if_type addr_if;
   data_if_type data_if;
   resp_if_type resp_if;
   rand int unsigned delay;
   axi_model#(T) slv_model;

   constraint delay_c {
      delay >= min_ready_delay;
      delay <= max_ready_delay;
   }

   axi_port_cfg cfg;

   function new(string name="axi_ready_driver", uvm_component parent=null);
      super.new(name, parent);
   endfunction // new

   `protect //begin protected region
   virtual function void build_phase(uvm_phase phase);
      super.build_phase(phase);
   endfunction // build_phase
   
   virtual function void connect_phase(uvm_phase phase);
      super.connect_phase(phase);
   endfunction // connect_phase

   task reset_phase(uvm_phase phase);
    //  phase.raise_objection(this);
    //  super.reset_phase(phase);
    //  if (channelType == AXI_ADDR) begin
    //     addr_if.dst_drv_cb.AxREADY <= '0;
    //     wait(addr_if.dst_drv_cb.resetn == 1'b1);
    //     repeat(10) @(addr_if.dst_drv_cb);
    //  end else if (channelType == AXI_DATA) begin
    //     data_if.dst_drv_cb.xREADY <= '0;
    //     wait(data_if.dst_drv_cb.resetn == 1'b1);
    //     repeat(10) @(data_if.dst_drv_cb);
    //  end else if (channelType == AXI_RESP) begin
    //     resp_if.dst_drv_cb.BREADY <= '0;
    //     wait(resp_if.dst_drv_cb.resetn == 1'b1);
    //     repeat(10) @(resp_if.dst_drv_cb);
    //  end
    //  `uvm_info(get_name(), "AXI_RESET_N deasserts", UVM_LOW)
    //  phase.drop_objection(this);
   endtask // reset_phase

   task reset_handler();
      if (channelType == AXI_ADDR) begin
         while (addr_if.dst_drv_cb.resetn === 1'b1 && (
               (cfg.unresponsive_slv_awready == 0 && direction == WRITE) ||
               (cfg.unresponsive_slv_arready == 0 && direction == READ))
         ) begin
            @(addr_if.dst_drv_cb);
         end
         addr_if.dst_drv_cb.AxREADY <= '0;
      end else if (channelType == AXI_DATA) begin
         while (data_if.dst_drv_cb.resetn === 1'b1) begin
            @(data_if.dst_drv_cb);
         end
         data_if.dst_drv_cb.xREADY <= '0;
      end else if (channelType == AXI_RESP) begin
         while (resp_if.dst_drv_cb.resetn === 1'b1) begin
            @(resp_if.dst_drv_cb);
         end
         resp_if.dst_drv_cb.BREADY <= '0;
      end
   endtask

   function void rand_delay();
      if (channelType == AXI_ADDR) begin
         min_ready_delay   = cfg.min_axready_delay;
         max_ready_delay   = cfg.max_axready_delay;
         ready_high_cycles = cfg.axready_high_cycles;
      end else if (channelType == AXI_DATA) begin
         min_ready_delay   = cfg.min_xready_delay;
         max_ready_delay   = cfg.max_xready_delay;
         ready_high_cycles = cfg.xready_high_cycles;
      end else if (channelType == AXI_RESP) begin
         min_ready_delay   = cfg.min_bready_delay;
         max_ready_delay   = cfg.max_bready_delay;
         ready_high_cycles = cfg.bready_high_cycles;
      end
      randomize(delay);
   endfunction

   task run_phase(uvm_phase phase);
      if (channelType == AXI_ADDR) begin
         addr_if.dst_drv_cb.AxREADY <= 1'b0;
         @(addr_if.dst_drv_cb);
         if (direction == WRITE) begin
            while (cfg.force_awready_low ==1) begin
               @(addr_if.dst_drv_cb);
            end
         end else if (direction == READ) begin
            while (cfg.force_arready_low ==1) begin
               @(addr_if.dst_drv_cb);
            end
         end
         min_ready_delay   = cfg.min_axready_delay;
         max_ready_delay   = cfg.max_axready_delay;
         ready_high_cycles = cfg.axready_high_cycles;
         repeat(cfg.initial_ready_delay_cycles) @(addr_if.dst_drv_cb);
      end else if (channelType == AXI_DATA) begin
         data_if.dst_drv_cb.xREADY <= 1'b0;
         @(data_if.dst_drv_cb);
         min_ready_delay   = cfg.min_xready_delay;
         max_ready_delay   = cfg.max_xready_delay;
         ready_high_cycles = cfg.xready_high_cycles;
         repeat(cfg.initial_ready_delay_cycles) @(data_if.dst_drv_cb);
      end else if (channelType == AXI_RESP) begin
         resp_if.dst_drv_cb.BREADY <= 1'b0;
         @(resp_if.dst_drv_cb);
         min_ready_delay   = cfg.min_bready_delay;
         max_ready_delay   = cfg.max_bready_delay;
         ready_high_cycles = cfg.bready_high_cycles;
         repeat(cfg.initial_ready_delay_cycles) @(resp_if.dst_drv_cb);
      end
      forever begin
         fork
            begin
               fork
                  reset_handler();
                  drive_if();
               join_any
            end
         join
         disable fork;
         if (channelType == AXI_ADDR) begin
            while (addr_if.src_drv_cb.resetn !== 1 || (
               (cfg.unresponsive_slv_awready == 1 && direction == WRITE) ||
               (cfg.unresponsive_slv_arready == 1 && direction == READ))
            ) begin
               @(addr_if.dst_drv_cb);
            end
         end else if (channelType == AXI_DATA) begin
            while (data_if.src_drv_cb.resetn !== 1) begin
               @(data_if.dst_drv_cb);
            end
         end else if (channelType == AXI_RESP) begin
            while (resp_if.src_drv_cb.resetn !== 1) begin
               @(resp_if.dst_drv_cb);
            end
         end
      end //forever
   endtask

   task drive_addr_using_delay();
      forever begin
         if ((cfg.unresponsive_slv_awready == 1 && direction == WRITE) || 
         (cfg.unresponsive_slv_arready == 1 && direction == READ)) begin
            addr_if.dst_drv_cb.AxREADY <= 1'b0;
            @(addr_if.dst_drv_cb);
         end  
         else if (addr_if.dst_drv_cb.resetn === 1'b1) begin
            if ((min_ready_delay == 0 && max_ready_delay == 0) || delay == 0) begin
               if (cfg.force_awready_low == 1) begin
                  addr_if.dst_drv_cb.AxREADY <= 1'b0;
               end else begin
                  addr_if.dst_drv_cb.AxREADY <= 1'b1;
               end
               @(addr_if.dst_drv_cb);
               while (addr_if.dst_drv_cb.AxVALID == 1'b0) begin
                  if (cfg.force_awready_low == 1) begin
                     addr_if.dst_drv_cb.AxREADY <= 1'b0;
                  end 
                  @(addr_if.dst_drv_cb);
               end
               rand_delay(); //randomize(delay); //next delay
            end else begin
               while (addr_if.dst_drv_cb.AxVALID == 1'b0) begin
                  if (cfg.force_awready_low == 1) begin
                     addr_if.dst_drv_cb.AxREADY <= 1'b0;
                  end 
                  @(addr_if.dst_drv_cb);
               end
               repeat(delay-1) @(addr_if.dst_drv_cb);
               if (cfg.force_awready_low == 1) begin
                  addr_if.dst_drv_cb.AxREADY <= 1'b0;
               end else begin
                  addr_if.dst_drv_cb.AxREADY <= 1'b1;
               end
               rand_delay(); //randomize(delay); //next delay
               @(addr_if.dst_drv_cb);
            end
            if (ready_high_cycles != 0) begin
               repeat(ready_high_cycles-1) @(addr_if.dst_drv_cb);
               addr_if.dst_drv_cb.AxREADY <= 1'b0;
               @(addr_if.dst_drv_cb);
            end
         end else begin
            addr_if.dst_drv_cb.AxREADY <= '0;
         end //if reset
      end //forever
   endtask

   task drive_addr_using_buffers();
      int unsigned buffer_size;
      int unsigned num_outstanding;

      if (direction == WRITE) begin
         buffer_size = cfg.slv_waddr_buffer_depth;
      end else begin
         buffer_size = cfg.slv_raddr_buffer_depth;
      end
      forever begin
         if ((cfg.unresponsive_slv_awready == 1 && direction == WRITE) ||
         (cfg.unresponsive_slv_arready == 1 && direction == READ) ) begin
            addr_if.dst_drv_cb.AxREADY <= 1'b0;
            @(addr_if.dst_drv_cb);
         end  
         else if (addr_if.dst_drv_cb.resetn === 1'b1) begin
            if (direction == WRITE) begin
               num_outstanding = slv_model.outstanding_wr_count; //get_num_pending_wr();
            end else begin
               num_outstanding = slv_model.outstanding_rd_count; //get_num_pending_rd();
            end
            if (num_outstanding < buffer_size) begin
               addr_if.dst_drv_cb.AxREADY <= 1'b1;
            end else begin
               addr_if.dst_drv_cb.AxREADY <= 1'b0;
            end
            @(addr_if.dst_drv_cb);
         end //if reset
      end //forever
   endtask

   task drive_if();
      //$display("%0t: %0s: drive_if :: %0s %0d %0d %0d", $time, get_full_name(), channelType.name(), min_ready_delay, max_ready_delay, ready_high_cycles);
      rand_delay();
      //randomize(delay); //initial delay
      if (channelType == AXI_ADDR) begin
         if (cfg.en_slv_buffers == 0) begin
            drive_addr_using_delay();
         end else begin
            drive_addr_using_buffers();
         end
      end else if (channelType == AXI_DATA) begin
         forever begin
            @(data_if.dst_drv_cb);
            if ((cfg.unresponsive_slv_wready == 1 && direction == WRITE) ||
            (cfg.unresponsive_mst_rready == 1 && direction == READ) ) begin
               data_if.dst_drv_cb.xREADY <= 1'b0;
            end
            else if (data_if.dst_drv_cb.resetn === 1'b1) begin
               if (!(min_ready_delay == 0 && max_ready_delay == 0)) begin
                  data_if.dst_drv_cb.xREADY <= 1'b0;
               end
               if (min_ready_delay == 0 && max_ready_delay == 0) begin
                  data_if.dst_drv_cb.xREADY <= 1'b1;
               end else begin
                  wait (data_if.dst_drv_cb.xVALID == 1'b1);
                  repeat(delay) @(data_if.dst_drv_cb);
                  data_if.dst_drv_cb.xREADY <= 1'b1;
                  rand_delay(); //randomize(delay); //next delay
               end
               if (ready_high_cycles != 0) begin
                  repeat(ready_high_cycles) @(data_if.dst_drv_cb);
                  data_if.dst_drv_cb.xREADY <= 1'b0;
               end
            end else begin
               data_if.dst_drv_cb.xREADY <= '0;
            end //if reset
         end //forever
      end else if (channelType == AXI_RESP) begin
         forever begin
            @(resp_if.dst_drv_cb);
            resp_if.dst_drv_cb.BREADY <= 1'b0;
            if (cfg.unresponsive_mst_bready == 1 && direction == WRITE) begin
               resp_if.dst_drv_cb.BREADY <= 1'b0;
            end else if (resp_if.dst_drv_cb.resetn === 1'b1) begin
               if (min_ready_delay == 0 && max_ready_delay == 0) begin
                  resp_if.dst_drv_cb.BREADY <= 1'b1;
               end else begin
                  wait (resp_if.dst_drv_cb.BVALID == 1'b1);
                  repeat(delay) @(resp_if.dst_drv_cb);
                  resp_if.dst_drv_cb.BREADY <= 1'b1;
                  rand_delay(); //randomize(delay); //next delay
               end
               if (ready_high_cycles != 0) begin
                  repeat(ready_high_cycles) @(resp_if.dst_drv_cb);
                  resp_if.dst_drv_cb.BREADY <= 1'b0;
               end
            end else begin
               resp_if.dst_drv_cb.BREADY <= '0;
            end //if reset
         end //forever
      end
   endtask

   `endprotect //end protected region

endclass
`endif
