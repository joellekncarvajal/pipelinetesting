/*
   ######################################################################################
 *      Signature IP Corporation Confidential and Proprietary Information               #
 *      Copyright 2022 Signature IP Corporation                                         #
 *      All Rights Reserved.                                                            #
 *      This is UNPUBLISHED PROPRIETARY SOURCE CODE OF Signature IP Corporation         #
 *      The copyright notice above does not evidence any actual or intended publication #
 *      of such source code.                                                            #
 * ######################################################################################

*/
`include "sig_test_base.sv"
`include "sig_axi_wr_rd_test.sv"
`include "sig_axi_burst_test.sv"
`include "sig_axi_mst_timing_test.sv"
`include "sig_axi_slv_timing_test.sv"
`include "sig_axi_write_interleaved_test.sv"
`include "sig_axi_read_interleaved_test.sv"
`include "sig_axi_error_response_test.sv"
